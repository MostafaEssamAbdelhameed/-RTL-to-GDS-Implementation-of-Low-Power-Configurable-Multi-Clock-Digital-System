module inv (
input q,
output d
);

assign d = !q ; 

endmodule 